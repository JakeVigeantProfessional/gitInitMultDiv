module bitwise_or(output_data,data1, data2);
input [31:0] data1, data2;
output [31:0] output_data;

or or0(output_data[0], data1[0], data2[0]);
or or1(output_data[1], data1[1], data2[1]);
or or2(output_data[2], data1[2], data2[2]);
or or3(output_data[3], data1[3], data2[3]);
or or4(output_data[4], data1[4], data2[4]);
or or5(output_data[5], data1[5], data2[5]);
or or6(output_data[6], data1[6], data2[6]);
or or7(output_data[7], data1[7], data2[7]);
or or8(output_data[8], data1[8], data2[8]);
or or9(output_data[9], data1[9], data2[9]);
or or10(output_data[10], data1[10], data2[10]);
or or11(output_data[11], data1[11], data2[11]);
or or12(output_data[12], data1[12], data2[12]);
or or13(output_data[13], data1[13], data2[13]);
or or14(output_data[14], data1[14], data2[14]);
or or15(output_data[15], data1[15], data2[15]);
or or16(output_data[16], data1[16], data2[16]);
or or17(output_data[17], data1[17], data2[17]);
or or18(output_data[18], data1[18], data2[18]);
or or19(output_data[19], data1[19], data2[19]);
or or20(output_data[20], data1[20], data2[20]);
or or21(output_data[21], data1[21], data2[21]);
or or22(output_data[22], data1[22], data2[22]);
or or23(output_data[23], data1[23], data2[23]);
or or24(output_data[24], data1[24], data2[24]);
or or25(output_data[25], data1[25], data2[25]);
or or26(output_data[26], data1[26], data2[26]);
or or27(output_data[27], data1[27], data2[27]);
or or28(output_data[28], data1[28], data2[28]);
or or29(output_data[29], data1[29], data2[29]);
or or30(output_data[30], data1[30], data2[30]);
or or31(output_data[31], data1[31], data2[31]);
endmodule